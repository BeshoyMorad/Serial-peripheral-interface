module MasterTB();

reg clk;
reg reset;
reg start;
reg [1:0] slaveSelect;
reg [7:0] masterDataToSend;
wire [7:0] masterDataReceived;
wire SCLK;
wire [0:2] CS;
wire MOSI;
reg MISO;

reg [7:0] data = 8'b01010011; // the data that will be sent to the master
reg [7:0] dataRecieved;  // the data recieved from the master
integer i;  // counter used to store data inside dataRecieved

Master M(
  clk, reset,
  start, slaveSelect, masterDataToSend, masterDataReceived,
  SCLK, CS, MOSI, MISO
);

initial 
begin
  clk = 1;
  reset = 1;
  #5 reset = 0;
  #15 start = 1;
  masterDataToSend = 8'b0010_0111;
  dataRecieved = 8'b0;
  slaveSelect = 0;
  #5 start = 0;

  // loop to send 8-bits to the master and get another 8-bits from it
  for(i=0 ; i<=7 ; i=i+1)
      begin
      if(i==0) begin
          MISO = data[0];
          #20 dataRecieved[0] = MOSI;
      end

      else begin
          #20 MISO = data[i];
          dataRecieved[i] = MOSI;
      end

      end

  #20;
  if(dataRecieved == masterDataToSend) 
      $display("From Master to Slave: Success");
  else 
      $display("From Master to Slave: Failure (Expected: %b, Received: %b)",  masterDataToSend, dataRecieved);
  if(masterDataReceived == data)
      $display("From Slave to Master: Success");
  else 
      $display("From Slave to Master: Failure (Expected: %b, Received: %b)", data, masterDataReceived);
  #10 $finish;

end

always #10 clk =~clk;

endmodule
